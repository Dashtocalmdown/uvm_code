program automatic test;
    import uvm_pkg::*;
    `include "uvm_macros.svh"
    //将之前的代码所创建的文件依次包含进来

    initial begin
        run_test();
    end

endprogram